// on_chip_with_keyboard_pio.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module on_chip_with_keyboard_pio (
		output wire [31:0] blue_export,            //            blue.export
		input  wire        clk_clk,                //             clk.clk
		output wire [31:0] exposure_export,        //        exposure.export
		output wire [31:0] green1_export,          //          green1.export
		output wire [31:0] green2_export,          //          green2.export
		output wire        mouse_click_export,     //     mouse_click.export
		output wire [11:0] mouse_x_export,         //         mouse_x.export
		output wire [11:0] mouse_y_export,         //         mouse_y.export
		output wire [1:0]  otg_hpi_address_export, // otg_hpi_address.export
		output wire        otg_hpi_cs_export,      //      otg_hpi_cs.export
		input  wire [15:0] otg_hpi_data_in_port,   //    otg_hpi_data.in_port
		output wire [15:0] otg_hpi_data_out_port,  //                .out_port
		output wire        otg_hpi_r_export,       //       otg_hpi_r.export
		output wire        otg_hpi_reset_export,   //   otg_hpi_reset.export
		output wire        otg_hpi_w_export,       //       otg_hpi_w.export
		output wire [31:0] red_export,             //             red.export
		input  wire        reset_reset_n           //           reset.reset_n
	);

	wire  [31:0] nios2_gen2_0_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                        // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [17:0] nios2_gen2_0_data_master_address;                            // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                         // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                               // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                              // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                          // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [17:0] nios2_gen2_0_instruction_master_address;                     // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                        // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;       // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;        // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;     // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;  // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [14:0] mm_interconnect_0_onchip_memory2_0_s1_address;               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_otg_hpi_address_s1_chipselect;             // mm_interconnect_0:otg_hpi_address_s1_chipselect -> otg_hpi_address:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_address_s1_readdata;               // otg_hpi_address:readdata -> mm_interconnect_0:otg_hpi_address_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_address_s1_address;                // mm_interconnect_0:otg_hpi_address_s1_address -> otg_hpi_address:address
	wire         mm_interconnect_0_otg_hpi_address_s1_write;                  // mm_interconnect_0:otg_hpi_address_s1_write -> otg_hpi_address:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_address_s1_writedata;              // mm_interconnect_0:otg_hpi_address_s1_writedata -> otg_hpi_address:writedata
	wire         mm_interconnect_0_otg_hpi_data_s1_chipselect;                // mm_interconnect_0:otg_hpi_data_s1_chipselect -> otg_hpi_data:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_data_s1_readdata;                  // otg_hpi_data:readdata -> mm_interconnect_0:otg_hpi_data_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_data_s1_address;                   // mm_interconnect_0:otg_hpi_data_s1_address -> otg_hpi_data:address
	wire         mm_interconnect_0_otg_hpi_data_s1_write;                     // mm_interconnect_0:otg_hpi_data_s1_write -> otg_hpi_data:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_data_s1_writedata;                 // mm_interconnect_0:otg_hpi_data_s1_writedata -> otg_hpi_data:writedata
	wire         mm_interconnect_0_otg_hpi_r_s1_chipselect;                   // mm_interconnect_0:otg_hpi_r_s1_chipselect -> otg_hpi_r:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_r_s1_readdata;                     // otg_hpi_r:readdata -> mm_interconnect_0:otg_hpi_r_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_r_s1_address;                      // mm_interconnect_0:otg_hpi_r_s1_address -> otg_hpi_r:address
	wire         mm_interconnect_0_otg_hpi_r_s1_write;                        // mm_interconnect_0:otg_hpi_r_s1_write -> otg_hpi_r:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_r_s1_writedata;                    // mm_interconnect_0:otg_hpi_r_s1_writedata -> otg_hpi_r:writedata
	wire         mm_interconnect_0_otg_hpi_w_s1_chipselect;                   // mm_interconnect_0:otg_hpi_w_s1_chipselect -> otg_hpi_w:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_w_s1_readdata;                     // otg_hpi_w:readdata -> mm_interconnect_0:otg_hpi_w_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_w_s1_address;                      // mm_interconnect_0:otg_hpi_w_s1_address -> otg_hpi_w:address
	wire         mm_interconnect_0_otg_hpi_w_s1_write;                        // mm_interconnect_0:otg_hpi_w_s1_write -> otg_hpi_w:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_w_s1_writedata;                    // mm_interconnect_0:otg_hpi_w_s1_writedata -> otg_hpi_w:writedata
	wire         mm_interconnect_0_otg_hpi_cs_s1_chipselect;                  // mm_interconnect_0:otg_hpi_cs_s1_chipselect -> otg_hpi_cs:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_cs_s1_readdata;                    // otg_hpi_cs:readdata -> mm_interconnect_0:otg_hpi_cs_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_cs_s1_address;                     // mm_interconnect_0:otg_hpi_cs_s1_address -> otg_hpi_cs:address
	wire         mm_interconnect_0_otg_hpi_cs_s1_write;                       // mm_interconnect_0:otg_hpi_cs_s1_write -> otg_hpi_cs:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_cs_s1_writedata;                   // mm_interconnect_0:otg_hpi_cs_s1_writedata -> otg_hpi_cs:writedata
	wire         mm_interconnect_0_otg_hpi_reset_s1_chipselect;               // mm_interconnect_0:otg_hpi_reset_s1_chipselect -> otg_hpi_reset:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_reset_s1_readdata;                 // otg_hpi_reset:readdata -> mm_interconnect_0:otg_hpi_reset_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_reset_s1_address;                  // mm_interconnect_0:otg_hpi_reset_s1_address -> otg_hpi_reset:address
	wire         mm_interconnect_0_otg_hpi_reset_s1_write;                    // mm_interconnect_0:otg_hpi_reset_s1_write -> otg_hpi_reset:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_reset_s1_writedata;                // mm_interconnect_0:otg_hpi_reset_s1_writedata -> otg_hpi_reset:writedata
	wire         mm_interconnect_0_mouse_x_s1_chipselect;                     // mm_interconnect_0:mouse_x_s1_chipselect -> mouse_x:chipselect
	wire  [31:0] mm_interconnect_0_mouse_x_s1_readdata;                       // mouse_x:readdata -> mm_interconnect_0:mouse_x_s1_readdata
	wire   [1:0] mm_interconnect_0_mouse_x_s1_address;                        // mm_interconnect_0:mouse_x_s1_address -> mouse_x:address
	wire         mm_interconnect_0_mouse_x_s1_write;                          // mm_interconnect_0:mouse_x_s1_write -> mouse_x:write_n
	wire  [31:0] mm_interconnect_0_mouse_x_s1_writedata;                      // mm_interconnect_0:mouse_x_s1_writedata -> mouse_x:writedata
	wire         mm_interconnect_0_mouse_y_s1_chipselect;                     // mm_interconnect_0:mouse_y_s1_chipselect -> mouse_y:chipselect
	wire  [31:0] mm_interconnect_0_mouse_y_s1_readdata;                       // mouse_y:readdata -> mm_interconnect_0:mouse_y_s1_readdata
	wire   [1:0] mm_interconnect_0_mouse_y_s1_address;                        // mm_interconnect_0:mouse_y_s1_address -> mouse_y:address
	wire         mm_interconnect_0_mouse_y_s1_write;                          // mm_interconnect_0:mouse_y_s1_write -> mouse_y:write_n
	wire  [31:0] mm_interconnect_0_mouse_y_s1_writedata;                      // mm_interconnect_0:mouse_y_s1_writedata -> mouse_y:writedata
	wire         mm_interconnect_0_mouse_click_s1_chipselect;                 // mm_interconnect_0:mouse_click_s1_chipselect -> mouse_click:chipselect
	wire  [31:0] mm_interconnect_0_mouse_click_s1_readdata;                   // mouse_click:readdata -> mm_interconnect_0:mouse_click_s1_readdata
	wire   [1:0] mm_interconnect_0_mouse_click_s1_address;                    // mm_interconnect_0:mouse_click_s1_address -> mouse_click:address
	wire         mm_interconnect_0_mouse_click_s1_write;                      // mm_interconnect_0:mouse_click_s1_write -> mouse_click:write_n
	wire  [31:0] mm_interconnect_0_mouse_click_s1_writedata;                  // mm_interconnect_0:mouse_click_s1_writedata -> mouse_click:writedata
	wire         mm_interconnect_0_exposure_s1_chipselect;                    // mm_interconnect_0:exposure_s1_chipselect -> exposure:chipselect
	wire  [31:0] mm_interconnect_0_exposure_s1_readdata;                      // exposure:readdata -> mm_interconnect_0:exposure_s1_readdata
	wire   [1:0] mm_interconnect_0_exposure_s1_address;                       // mm_interconnect_0:exposure_s1_address -> exposure:address
	wire         mm_interconnect_0_exposure_s1_write;                         // mm_interconnect_0:exposure_s1_write -> exposure:write_n
	wire  [31:0] mm_interconnect_0_exposure_s1_writedata;                     // mm_interconnect_0:exposure_s1_writedata -> exposure:writedata
	wire         mm_interconnect_0_green1_s1_chipselect;                      // mm_interconnect_0:green1_s1_chipselect -> green1:chipselect
	wire  [31:0] mm_interconnect_0_green1_s1_readdata;                        // green1:readdata -> mm_interconnect_0:green1_s1_readdata
	wire   [1:0] mm_interconnect_0_green1_s1_address;                         // mm_interconnect_0:green1_s1_address -> green1:address
	wire         mm_interconnect_0_green1_s1_write;                           // mm_interconnect_0:green1_s1_write -> green1:write_n
	wire  [31:0] mm_interconnect_0_green1_s1_writedata;                       // mm_interconnect_0:green1_s1_writedata -> green1:writedata
	wire         mm_interconnect_0_green2_s1_chipselect;                      // mm_interconnect_0:green2_s1_chipselect -> green2:chipselect
	wire  [31:0] mm_interconnect_0_green2_s1_readdata;                        // green2:readdata -> mm_interconnect_0:green2_s1_readdata
	wire   [1:0] mm_interconnect_0_green2_s1_address;                         // mm_interconnect_0:green2_s1_address -> green2:address
	wire         mm_interconnect_0_green2_s1_write;                           // mm_interconnect_0:green2_s1_write -> green2:write_n
	wire  [31:0] mm_interconnect_0_green2_s1_writedata;                       // mm_interconnect_0:green2_s1_writedata -> green2:writedata
	wire         mm_interconnect_0_red_s1_chipselect;                         // mm_interconnect_0:red_s1_chipselect -> red:chipselect
	wire  [31:0] mm_interconnect_0_red_s1_readdata;                           // red:readdata -> mm_interconnect_0:red_s1_readdata
	wire   [1:0] mm_interconnect_0_red_s1_address;                            // mm_interconnect_0:red_s1_address -> red:address
	wire         mm_interconnect_0_red_s1_write;                              // mm_interconnect_0:red_s1_write -> red:write_n
	wire  [31:0] mm_interconnect_0_red_s1_writedata;                          // mm_interconnect_0:red_s1_writedata -> red:writedata
	wire         mm_interconnect_0_blue_s1_chipselect;                        // mm_interconnect_0:blue_s1_chipselect -> blue:chipselect
	wire  [31:0] mm_interconnect_0_blue_s1_readdata;                          // blue:readdata -> mm_interconnect_0:blue_s1_readdata
	wire   [1:0] mm_interconnect_0_blue_s1_address;                           // mm_interconnect_0:blue_s1_address -> blue:address
	wire         mm_interconnect_0_blue_s1_write;                             // mm_interconnect_0:blue_s1_write -> blue:write_n
	wire  [31:0] mm_interconnect_0_blue_s1_writedata;                         // mm_interconnect_0:blue_s1_writedata -> blue:writedata
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [blue:reset_n, exposure:reset_n, green1:reset_n, green2:reset_n, jtag_uart_0:rst_n, mm_interconnect_0:jtag_uart_0_reset_reset_bridge_in_reset_reset, mouse_click:reset_n, mouse_x:reset_n, mouse_y:reset_n, onchip_memory2_0:reset, otg_hpi_address:reset_n, otg_hpi_cs:reset_n, otg_hpi_data:reset_n, otg_hpi_r:reset_n, otg_hpi_reset:reset_n, otg_hpi_w:reset_n, red:reset_n, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, rst_translator_001:in_reset, sysid_qsys_0:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                      // rst_controller_001:reset_req -> [nios2_gen2_0:reset_req, rst_translator_001:reset_req_in]
	wire         nios2_gen2_0_debug_reset_request_reset;                      // nios2_gen2_0:debug_reset_request -> rst_controller_001:reset_in1

	on_chip_with_keyboard_pio_blue blue (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_blue_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_blue_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_blue_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_blue_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_blue_s1_readdata),   //                    .readdata
		.out_port   (blue_export)                           // external_connection.export
	);

	on_chip_with_keyboard_pio_blue exposure (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_exposure_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_exposure_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_exposure_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_exposure_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_exposure_s1_readdata),   //                    .readdata
		.out_port   (exposure_export)                           // external_connection.export
	);

	on_chip_with_keyboard_pio_blue green1 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_green1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_green1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_green1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_green1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_green1_s1_readdata),   //                    .readdata
		.out_port   (green1_export)                           // external_connection.export
	);

	on_chip_with_keyboard_pio_blue green2 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_green2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_green2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_green2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_green2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_green2_s1_readdata),   //                    .readdata
		.out_port   (green2_export)                           // external_connection.export
	);

	on_chip_with_keyboard_pio_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	on_chip_with_keyboard_pio_mouse_click mouse_click (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_mouse_click_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_mouse_click_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_mouse_click_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_mouse_click_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_mouse_click_s1_readdata),   //                    .readdata
		.out_port   (mouse_click_export)                           // external_connection.export
	);

	on_chip_with_keyboard_pio_mouse_x mouse_x (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_mouse_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_mouse_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_mouse_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_mouse_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_mouse_x_s1_readdata),   //                    .readdata
		.out_port   (mouse_x_export)                           // external_connection.export
	);

	on_chip_with_keyboard_pio_mouse_x mouse_y (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_mouse_y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_mouse_y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_mouse_y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_mouse_y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_mouse_y_s1_readdata),   //                    .readdata
		.out_port   (mouse_y_export)                           // external_connection.export
	);

	on_chip_with_keyboard_pio_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	on_chip_with_keyboard_pio_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	on_chip_with_keyboard_pio_otg_hpi_address otg_hpi_address (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_address_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_address_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_address_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_address_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_address_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_address_export)                           // external_connection.export
	);

	on_chip_with_keyboard_pio_mouse_click otg_hpi_cs (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_cs_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_cs_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_cs_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_cs_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_cs_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_cs_export)                           // external_connection.export
	);

	on_chip_with_keyboard_pio_otg_hpi_data otg_hpi_data (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_data_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_data_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_data_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_data_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_data_s1_readdata),   //                    .readdata
		.in_port    (otg_hpi_data_in_port),                         // external_connection.export
		.out_port   (otg_hpi_data_out_port)                         //                    .export
	);

	on_chip_with_keyboard_pio_mouse_click otg_hpi_r (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_r_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_r_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_r_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_r_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_r_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_r_export)                           // external_connection.export
	);

	on_chip_with_keyboard_pio_mouse_click otg_hpi_reset (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_reset_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_reset_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_reset_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_reset_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_reset_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_reset_export)                           // external_connection.export
	);

	on_chip_with_keyboard_pio_mouse_click otg_hpi_w (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_w_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_w_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_w_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_w_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_w_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_w_export)                           // external_connection.export
	);

	on_chip_with_keyboard_pio_blue red (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_red_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_red_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_red_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_red_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_red_s1_readdata),   //                    .readdata
		.out_port   (red_export)                           // external_connection.export
	);

	on_chip_with_keyboard_pio_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	on_chip_with_keyboard_pio_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                     //                                clk_0_clk.clk
		.jtag_uart_0_reset_reset_bridge_in_reset_reset  (rst_controller_reset_out_reset),                              //  jtag_uart_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                            //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                        //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                         //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                               //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                           //                                         .readdata
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                              //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                          //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                        //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                     //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                 //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                        //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                    //                                         .readdata
		.blue_s1_address                                (mm_interconnect_0_blue_s1_address),                           //                                  blue_s1.address
		.blue_s1_write                                  (mm_interconnect_0_blue_s1_write),                             //                                         .write
		.blue_s1_readdata                               (mm_interconnect_0_blue_s1_readdata),                          //                                         .readdata
		.blue_s1_writedata                              (mm_interconnect_0_blue_s1_writedata),                         //                                         .writedata
		.blue_s1_chipselect                             (mm_interconnect_0_blue_s1_chipselect),                        //                                         .chipselect
		.exposure_s1_address                            (mm_interconnect_0_exposure_s1_address),                       //                              exposure_s1.address
		.exposure_s1_write                              (mm_interconnect_0_exposure_s1_write),                         //                                         .write
		.exposure_s1_readdata                           (mm_interconnect_0_exposure_s1_readdata),                      //                                         .readdata
		.exposure_s1_writedata                          (mm_interconnect_0_exposure_s1_writedata),                     //                                         .writedata
		.exposure_s1_chipselect                         (mm_interconnect_0_exposure_s1_chipselect),                    //                                         .chipselect
		.green1_s1_address                              (mm_interconnect_0_green1_s1_address),                         //                                green1_s1.address
		.green1_s1_write                                (mm_interconnect_0_green1_s1_write),                           //                                         .write
		.green1_s1_readdata                             (mm_interconnect_0_green1_s1_readdata),                        //                                         .readdata
		.green1_s1_writedata                            (mm_interconnect_0_green1_s1_writedata),                       //                                         .writedata
		.green1_s1_chipselect                           (mm_interconnect_0_green1_s1_chipselect),                      //                                         .chipselect
		.green2_s1_address                              (mm_interconnect_0_green2_s1_address),                         //                                green2_s1.address
		.green2_s1_write                                (mm_interconnect_0_green2_s1_write),                           //                                         .write
		.green2_s1_readdata                             (mm_interconnect_0_green2_s1_readdata),                        //                                         .readdata
		.green2_s1_writedata                            (mm_interconnect_0_green2_s1_writedata),                       //                                         .writedata
		.green2_s1_chipselect                           (mm_interconnect_0_green2_s1_chipselect),                      //                                         .chipselect
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.mouse_click_s1_address                         (mm_interconnect_0_mouse_click_s1_address),                    //                           mouse_click_s1.address
		.mouse_click_s1_write                           (mm_interconnect_0_mouse_click_s1_write),                      //                                         .write
		.mouse_click_s1_readdata                        (mm_interconnect_0_mouse_click_s1_readdata),                   //                                         .readdata
		.mouse_click_s1_writedata                       (mm_interconnect_0_mouse_click_s1_writedata),                  //                                         .writedata
		.mouse_click_s1_chipselect                      (mm_interconnect_0_mouse_click_s1_chipselect),                 //                                         .chipselect
		.mouse_x_s1_address                             (mm_interconnect_0_mouse_x_s1_address),                        //                               mouse_x_s1.address
		.mouse_x_s1_write                               (mm_interconnect_0_mouse_x_s1_write),                          //                                         .write
		.mouse_x_s1_readdata                            (mm_interconnect_0_mouse_x_s1_readdata),                       //                                         .readdata
		.mouse_x_s1_writedata                           (mm_interconnect_0_mouse_x_s1_writedata),                      //                                         .writedata
		.mouse_x_s1_chipselect                          (mm_interconnect_0_mouse_x_s1_chipselect),                     //                                         .chipselect
		.mouse_y_s1_address                             (mm_interconnect_0_mouse_y_s1_address),                        //                               mouse_y_s1.address
		.mouse_y_s1_write                               (mm_interconnect_0_mouse_y_s1_write),                          //                                         .write
		.mouse_y_s1_readdata                            (mm_interconnect_0_mouse_y_s1_readdata),                       //                                         .readdata
		.mouse_y_s1_writedata                           (mm_interconnect_0_mouse_y_s1_writedata),                      //                                         .writedata
		.mouse_y_s1_chipselect                          (mm_interconnect_0_mouse_y_s1_chipselect),                     //                                         .chipselect
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),      //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),        //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),         //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),     //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),    //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),   //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),  //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),  //                                         .debugaccess
		.onchip_memory2_0_s1_address                    (mm_interconnect_0_onchip_memory2_0_s1_address),               //                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                      (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                         .write
		.onchip_memory2_0_s1_readdata                   (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                         .readdata
		.onchip_memory2_0_s1_writedata                  (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                         .writedata
		.onchip_memory2_0_s1_byteenable                 (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                         .byteenable
		.onchip_memory2_0_s1_chipselect                 (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                         .chipselect
		.onchip_memory2_0_s1_clken                      (mm_interconnect_0_onchip_memory2_0_s1_clken),                 //                                         .clken
		.otg_hpi_address_s1_address                     (mm_interconnect_0_otg_hpi_address_s1_address),                //                       otg_hpi_address_s1.address
		.otg_hpi_address_s1_write                       (mm_interconnect_0_otg_hpi_address_s1_write),                  //                                         .write
		.otg_hpi_address_s1_readdata                    (mm_interconnect_0_otg_hpi_address_s1_readdata),               //                                         .readdata
		.otg_hpi_address_s1_writedata                   (mm_interconnect_0_otg_hpi_address_s1_writedata),              //                                         .writedata
		.otg_hpi_address_s1_chipselect                  (mm_interconnect_0_otg_hpi_address_s1_chipselect),             //                                         .chipselect
		.otg_hpi_cs_s1_address                          (mm_interconnect_0_otg_hpi_cs_s1_address),                     //                            otg_hpi_cs_s1.address
		.otg_hpi_cs_s1_write                            (mm_interconnect_0_otg_hpi_cs_s1_write),                       //                                         .write
		.otg_hpi_cs_s1_readdata                         (mm_interconnect_0_otg_hpi_cs_s1_readdata),                    //                                         .readdata
		.otg_hpi_cs_s1_writedata                        (mm_interconnect_0_otg_hpi_cs_s1_writedata),                   //                                         .writedata
		.otg_hpi_cs_s1_chipselect                       (mm_interconnect_0_otg_hpi_cs_s1_chipselect),                  //                                         .chipselect
		.otg_hpi_data_s1_address                        (mm_interconnect_0_otg_hpi_data_s1_address),                   //                          otg_hpi_data_s1.address
		.otg_hpi_data_s1_write                          (mm_interconnect_0_otg_hpi_data_s1_write),                     //                                         .write
		.otg_hpi_data_s1_readdata                       (mm_interconnect_0_otg_hpi_data_s1_readdata),                  //                                         .readdata
		.otg_hpi_data_s1_writedata                      (mm_interconnect_0_otg_hpi_data_s1_writedata),                 //                                         .writedata
		.otg_hpi_data_s1_chipselect                     (mm_interconnect_0_otg_hpi_data_s1_chipselect),                //                                         .chipselect
		.otg_hpi_r_s1_address                           (mm_interconnect_0_otg_hpi_r_s1_address),                      //                             otg_hpi_r_s1.address
		.otg_hpi_r_s1_write                             (mm_interconnect_0_otg_hpi_r_s1_write),                        //                                         .write
		.otg_hpi_r_s1_readdata                          (mm_interconnect_0_otg_hpi_r_s1_readdata),                     //                                         .readdata
		.otg_hpi_r_s1_writedata                         (mm_interconnect_0_otg_hpi_r_s1_writedata),                    //                                         .writedata
		.otg_hpi_r_s1_chipselect                        (mm_interconnect_0_otg_hpi_r_s1_chipselect),                   //                                         .chipselect
		.otg_hpi_reset_s1_address                       (mm_interconnect_0_otg_hpi_reset_s1_address),                  //                         otg_hpi_reset_s1.address
		.otg_hpi_reset_s1_write                         (mm_interconnect_0_otg_hpi_reset_s1_write),                    //                                         .write
		.otg_hpi_reset_s1_readdata                      (mm_interconnect_0_otg_hpi_reset_s1_readdata),                 //                                         .readdata
		.otg_hpi_reset_s1_writedata                     (mm_interconnect_0_otg_hpi_reset_s1_writedata),                //                                         .writedata
		.otg_hpi_reset_s1_chipselect                    (mm_interconnect_0_otg_hpi_reset_s1_chipselect),               //                                         .chipselect
		.otg_hpi_w_s1_address                           (mm_interconnect_0_otg_hpi_w_s1_address),                      //                             otg_hpi_w_s1.address
		.otg_hpi_w_s1_write                             (mm_interconnect_0_otg_hpi_w_s1_write),                        //                                         .write
		.otg_hpi_w_s1_readdata                          (mm_interconnect_0_otg_hpi_w_s1_readdata),                     //                                         .readdata
		.otg_hpi_w_s1_writedata                         (mm_interconnect_0_otg_hpi_w_s1_writedata),                    //                                         .writedata
		.otg_hpi_w_s1_chipselect                        (mm_interconnect_0_otg_hpi_w_s1_chipselect),                   //                                         .chipselect
		.red_s1_address                                 (mm_interconnect_0_red_s1_address),                            //                                   red_s1.address
		.red_s1_write                                   (mm_interconnect_0_red_s1_write),                              //                                         .write
		.red_s1_readdata                                (mm_interconnect_0_red_s1_readdata),                           //                                         .readdata
		.red_s1_writedata                               (mm_interconnect_0_red_s1_writedata),                          //                                         .writedata
		.red_s1_chipselect                              (mm_interconnect_0_red_s1_chipselect),                         //                                         .chipselect
		.sysid_qsys_0_control_slave_address             (mm_interconnect_0_sysid_qsys_0_control_slave_address),        //               sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata            (mm_interconnect_0_sysid_qsys_0_control_slave_readdata)        //                                         .readdata
	);

	on_chip_with_keyboard_pio_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.sender_irq    (nios2_gen2_0_irq_irq)                //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
